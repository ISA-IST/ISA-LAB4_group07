
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY dadda_tree IS
PORT (
	pp0, pp1, pp2, pp3, pp4, pp5, pp6, pp7, pp8, pp9, 
	pp10, pp11, pp12, pp13, pp14, pp15: IN STD_LOGIC_VECTOR(32 downto 0);
	pp16: IN STD_LOGIC_VECTOR(31 downto 0);
	s: IN STD_LOGIC_VECTOR(15 downto 0);
	s_n: IN STD_LOGIC_VECTOR(15 downto 0);
	addend1_out, addend2_out: OUT STD_LOGIC_VECTOR(62 downto 0);
	M_lsb: OUT STD_LOGIC
);
END dadda_tree;

ARCHITECTURE struct OF dadda_tree IS

	COMPONENT FA IS
	PORT(
		a, b, c_in : IN std_logic;
		s, c_out : OUT std_logic);
	END COMPONENT;

	COMPONENT HA IS
	PORT(
		a, b : IN std_logic;
		s, c_out : OUT std_logic);
	END COMPONENT;

	SIGNAL sum_0, c_out_0: STD_LOGIC_VECTOR (51 downto 0);
	SIGNAL sum_1, c_out_1: STD_LOGIC_VECTOR (115 downto 0);
	SIGNAL sum_2, c_out_2: STD_LOGIC_VECTOR (128 downto 0);
	SIGNAL sum_3, c_out_3: STD_LOGIC_VECTOR (105 downto 0);
	SIGNAL sum_4, c_out_4: STD_LOGIC_VECTOR (58 downto 0);
	SIGNAL sum_5, c_out_5: STD_LOGIC_VECTOR (61 downto 0);
	SIGNAL sum_6, c_out_6: STD_LOGIC;

BEGIN

	HA_0_0 : HA port map (A=>pp12(0), B=>s(12), S=>sum_0(0) , C_out=>c_out_0(0));
	HA_0_1 : HA port map (A=>pp11(3), B=>pp12(1), S=>sum_0(1) , C_out=>c_out_0(1));
	FA_0_2 : FA port map (A=>pp12(2), B=>pp13(0), C_in=>s(13), S=>sum_0(2) , C_out=>c_out_0(2));
	HA_0_3 : HA port map (A=>pp10(6), B=>pp11(4), S=>sum_0(3) , C_out=>c_out_0(3));
	FA_0_4 : FA port map (A=>pp11(5), B=>pp12(3), C_in=>pp13(1), S=>sum_0(4) , C_out=>c_out_0(4));
	HA_0_5 : HA port map (A=>pp9(9), B=>pp10(7), S=>sum_0(5) , C_out=>c_out_0(5));
	FA_0_6 : FA port map (A=>pp13(2), B=>pp14(0), C_in=>s(14), S=>sum_0(6) , C_out=>c_out_0(6));
	FA_0_7 : FA port map (A=>pp10(8), B=>pp11(6), C_in=>pp12(4), S=>sum_0(7) , C_out=>c_out_0(7));
	HA_0_8 : HA port map (A=>pp8(12), B=>pp9(10), S=>sum_0(8) , C_out=>c_out_0(8));
	FA_0_9 : FA port map (A=>pp12(5), B=>pp13(3), C_in=>pp14(1), S=>sum_0(9) , C_out=>c_out_0(9));
	FA_0_10 : FA port map (A=>pp9(11), B=>pp10(9), C_in=>pp11(7), S=>sum_0(10) , C_out=>c_out_0(10));
	HA_0_11 : HA port map (A=>pp7(15), B=>pp8(13), S=>sum_0(11) , C_out=>c_out_0(11));
	FA_0_12 : FA port map (A=>pp14(2), B=>pp15(0), C_in=>s(15), S=>sum_0(12) , C_out=>c_out_0(12));
	FA_0_13 : FA port map (A=>pp11(8), B=>pp12(6), C_in=>pp13(4), S=>sum_0(13) , C_out=>c_out_0(13));
	FA_0_14 : FA port map (A=>pp8(14), B=>pp9(12), C_in=>pp10(10), S=>sum_0(14) , C_out=>c_out_0(14));
	HA_0_15 : HA port map (A=>pp6(18), B=>pp7(16), S=>sum_0(15) , C_out=>c_out_0(15));
	FA_0_16 : FA port map (A=>pp13(5), B=>pp14(3), C_in=>pp15(1), S=>sum_0(16) , C_out=>c_out_0(16));
	FA_0_17 : FA port map (A=>pp10(11), B=>pp11(9), C_in=>pp12(7), S=>sum_0(17) , C_out=>c_out_0(17));
	FA_0_18 : FA port map (A=>pp7(17), B=>pp8(15), C_in=>pp9(13), S=>sum_0(18) , C_out=>c_out_0(18));
	HA_0_19 : HA port map (A=>pp5(21), B=>pp6(19), S=>sum_0(19) , C_out=>c_out_0(19));
	FA_0_20 : FA port map (A=>pp14(4), B=>pp15(2), C_in=>pp16(0), S=>sum_0(20) , C_out=>c_out_0(20));
	FA_0_21 : FA port map (A=>pp11(10), B=>pp12(8), C_in=>pp13(6), S=>sum_0(21) , C_out=>c_out_0(21));
	FA_0_22 : FA port map (A=>pp8(16), B=>pp9(14), C_in=>pp10(12), S=>sum_0(22) , C_out=>c_out_0(22));
	FA_0_23 : FA port map (A=>pp5(22), B=>pp6(20), C_in=>pp7(18), S=>sum_0(23) , C_out=>c_out_0(23));
	FA_0_24 : FA port map (A=>pp14(5), B=>pp15(3), C_in=>pp16(1), S=>sum_0(24) , C_out=>c_out_0(24));
	FA_0_25 : FA port map (A=>pp11(11), B=>pp12(9), C_in=>pp13(7), S=>sum_0(25) , C_out=>c_out_0(25));
	FA_0_26 : FA port map (A=>pp8(17), B=>pp9(15), C_in=>pp10(13), S=>sum_0(26) , C_out=>c_out_0(26));
	FA_0_27 : FA port map (A=>pp5(23), B=>pp6(21), C_in=>pp7(19), S=>sum_0(27) , C_out=>c_out_0(27));
	FA_0_28 : FA port map (A=>pp14(6), B=>pp15(4), C_in=>pp16(2), S=>sum_0(28) , C_out=>c_out_0(28));
	FA_0_29 : FA port map (A=>pp11(12), B=>pp12(10), C_in=>pp13(8), S=>sum_0(29) , C_out=>c_out_0(29));
	FA_0_30 : FA port map (A=>pp8(18), B=>pp9(16), C_in=>pp10(14), S=>sum_0(30) , C_out=>c_out_0(30));
	FA_0_31 : FA port map (A=>pp5(24), B=>pp6(22), C_in=>pp7(20), S=>sum_0(31) , C_out=>c_out_0(31));
	FA_0_32 : FA port map (A=>pp14(7), B=>pp15(5), C_in=>pp16(3), S=>sum_0(32) , C_out=>c_out_0(32));
	FA_0_33 : FA port map (A=>pp11(13), B=>pp12(11), C_in=>pp13(9), S=>sum_0(33) , C_out=>c_out_0(33));
	FA_0_34 : FA port map (A=>pp8(19), B=>pp9(17), C_in=>pp10(15), S=>sum_0(34) , C_out=>c_out_0(34));
	FA_0_35 : FA port map (A=>pp5(25), B=>pp6(23), C_in=>pp7(21), S=>sum_0(35) , C_out=>c_out_0(35));
	FA_0_36 : FA port map (A=>pp14(8), B=>pp15(6), C_in=>pp16(4), S=>sum_0(36) , C_out=>c_out_0(36));
	FA_0_37 : FA port map (A=>pp11(14), B=>pp12(12), C_in=>pp13(10), S=>sum_0(37) , C_out=>c_out_0(37));
	FA_0_38 : FA port map (A=>pp8(20), B=>pp9(18), C_in=>pp10(16), S=>sum_0(38) , C_out=>c_out_0(38));
	HA_0_39 : HA port map (A=>pp6(24), B=>pp7(22), S=>sum_0(39) , C_out=>c_out_0(39));
	FA_0_40 : FA port map (A=>pp14(9), B=>pp15(7), C_in=>pp16(5), S=>sum_0(40) , C_out=>c_out_0(40));
	FA_0_41 : FA port map (A=>pp11(15), B=>pp12(13), C_in=>pp13(11), S=>sum_0(41) , C_out=>c_out_0(41));
	FA_0_42 : FA port map (A=>pp8(21), B=>pp9(19), C_in=>pp10(17), S=>sum_0(42) , C_out=>c_out_0(42));
	FA_0_43 : FA port map (A=>pp14(10), B=>pp15(8), C_in=>pp16(6), S=>sum_0(43) , C_out=>c_out_0(43));
	FA_0_44 : FA port map (A=>pp11(16), B=>pp12(14), C_in=>pp13(12), S=>sum_0(44) , C_out=>c_out_0(44));
	HA_0_45 : HA port map (A=>pp9(20), B=>pp10(18), S=>sum_0(45) , C_out=>c_out_0(45));
	FA_0_46 : FA port map (A=>pp14(11), B=>pp15(9), C_in=>pp16(7), S=>sum_0(46) , C_out=>c_out_0(46));
	FA_0_47 : FA port map (A=>pp11(17), B=>pp12(15), C_in=>pp13(13), S=>sum_0(47) , C_out=>c_out_0(47));
	FA_0_48 : FA port map (A=>pp14(12), B=>pp15(10), C_in=>pp16(8), S=>sum_0(48) , C_out=>c_out_0(48));
	HA_0_49 : HA port map (A=>pp12(16), B=>pp13(14), S=>sum_0(49) , C_out=>c_out_0(49));
	FA_0_50 : FA port map (A=>pp14(13), B=>pp15(11), C_in=>pp16(9), S=>sum_0(50) , C_out=>c_out_0(50));
	HA_0_51 : HA port map (A=>pp15(12), B=>pp16(10), S=>sum_0(51) , C_out=>c_out_0(51));
	HA_1_0 : HA port map (A=>pp8(0), B=>s(8), S=>sum_1(0) , C_out=>c_out_1(0));
	HA_1_1 : HA port map (A=>pp7(3), B=>pp8(1), S=>sum_1(1) , C_out=>c_out_1(1));
	FA_1_2 : FA port map (A=>pp8(2), B=>pp9(0), C_in=>s(9), S=>sum_1(2) , C_out=>c_out_1(2));
	HA_1_3 : HA port map (A=>pp6(6), B=>pp7(4), S=>sum_1(3) , C_out=>c_out_1(3));
	FA_1_4 : FA port map (A=>pp7(5), B=>pp8(3), C_in=>pp9(1), S=>sum_1(4) , C_out=>c_out_1(4));
	HA_1_5 : HA port map (A=>pp5(9), B=>pp6(7), S=>sum_1(5) , C_out=>c_out_1(5));
	FA_1_6 : FA port map (A=>pp9(2), B=>pp10(0), C_in=>s(10), S=>sum_1(6) , C_out=>c_out_1(6));
	FA_1_7 : FA port map (A=>pp6(8), B=>pp7(6), C_in=>pp8(4), S=>sum_1(7) , C_out=>c_out_1(7));
	HA_1_8 : HA port map (A=>pp4(12), B=>pp5(10), S=>sum_1(8) , C_out=>c_out_1(8));
	FA_1_9 : FA port map (A=>pp8(5), B=>pp9(3), C_in=>pp10(1), S=>sum_1(9) , C_out=>c_out_1(9));
	FA_1_10 : FA port map (A=>pp5(11), B=>pp6(9), C_in=>pp7(7), S=>sum_1(10) , C_out=>c_out_1(10));
	HA_1_11 : HA port map (A=>pp3(15), B=>pp4(13), S=>sum_1(11) , C_out=>c_out_1(11));
	FA_1_12 : FA port map (A=>pp10(2), B=>pp11(0), C_in=>s(11), S=>sum_1(12) , C_out=>c_out_1(12));
	FA_1_13 : FA port map (A=>pp7(8), B=>pp8(6), C_in=>pp9(4), S=>sum_1(13) , C_out=>c_out_1(13));
	FA_1_14 : FA port map (A=>pp4(14), B=>pp5(12), C_in=>pp6(10), S=>sum_1(14) , C_out=>c_out_1(14));
	HA_1_15 : HA port map (A=>pp2(18), B=>pp3(16), S=>sum_1(15) , C_out=>c_out_1(15));
	FA_1_16 : FA port map (A=>pp9(5), B=>pp10(3), C_in=>pp11(1), S=>sum_1(16) , C_out=>c_out_1(16));
	FA_1_17 : FA port map (A=>pp6(11), B=>pp7(9), C_in=>pp8(7), S=>sum_1(17) , C_out=>c_out_1(17));
	FA_1_18 : FA port map (A=>pp3(17), B=>pp4(15), C_in=>pp5(13), S=>sum_1(18) , C_out=>c_out_1(18));
	HA_1_19 : HA port map (A=>pp1(21), B=>pp2(19), S=>sum_1(19) , C_out=>c_out_1(19));
	FA_1_20 : FA port map (A=>pp9(6), B=>pp10(4), C_in=>pp11(2), S=>sum_1(20) , C_out=>c_out_1(20));
	FA_1_21 : FA port map (A=>pp6(12), B=>pp7(10), C_in=>pp8(8), S=>sum_1(21) , C_out=>c_out_1(21));
	FA_1_22 : FA port map (A=>pp3(18), B=>pp4(16), C_in=>pp5(14), S=>sum_1(22) , C_out=>c_out_1(22));
	FA_1_23 : FA port map (A=>pp0(24), B=>pp1(22), C_in=>pp2(20), S=>sum_1(23) , C_out=>c_out_1(23));
	FA_1_24 : FA port map (A=>pp8(9), B=>pp9(7), C_in=>pp10(5), S=>sum_1(24) , C_out=>c_out_1(24));
	FA_1_25 : FA port map (A=>pp5(15), B=>pp6(13), C_in=>pp7(11), S=>sum_1(25) , C_out=>c_out_1(25));
	FA_1_26 : FA port map (A=>pp2(21), B=>pp3(19), C_in=>pp4(17), S=>sum_1(26) , C_out=>c_out_1(26));
	FA_1_27 : FA port map (A=>c_out_0(0), B=>pp0(25), C_in=>pp1(23), S=>sum_1(27) , C_out=>c_out_1(27));
	FA_1_28 : FA port map (A=>pp7(12), B=>pp8(10), C_in=>pp9(8), S=>sum_1(28) , C_out=>c_out_1(28));
	FA_1_29 : FA port map (A=>pp4(18), B=>pp5(16), C_in=>pp6(14), S=>sum_1(29) , C_out=>c_out_1(29));
	FA_1_30 : FA port map (A=>pp1(24), B=>pp2(22), C_in=>pp3(20), S=>sum_1(30) , C_out=>c_out_1(30));
	FA_1_31 : FA port map (A=>sum_0(2), B=>c_out_0(1), C_in=>pp0(26), S=>sum_1(31) , C_out=>c_out_1(31));
	FA_1_32 : FA port map (A=>pp6(15), B=>pp7(13), C_in=>pp8(11), S=>sum_1(32) , C_out=>c_out_1(32));
	FA_1_33 : FA port map (A=>pp3(21), B=>pp4(19), C_in=>pp5(17), S=>sum_1(33) , C_out=>c_out_1(33));
	FA_1_34 : FA port map (A=>pp0(27), B=>pp1(25), C_in=>pp2(23), S=>sum_1(34) , C_out=>c_out_1(34));
	FA_1_35 : FA port map (A=>sum_0(4), B=>c_out_0(3), C_in=>c_out_0(2), S=>sum_1(35) , C_out=>c_out_1(35));
	FA_1_36 : FA port map (A=>pp5(18), B=>pp6(16), C_in=>pp7(14), S=>sum_1(36) , C_out=>c_out_1(36));
	FA_1_37 : FA port map (A=>pp2(24), B=>pp3(22), C_in=>pp4(20), S=>sum_1(37) , C_out=>c_out_1(37));
	FA_1_38 : FA port map (A=>c_out_0(4), B=>pp0(28), C_in=>pp1(26), S=>sum_1(38) , C_out=>c_out_1(38));
	FA_1_39 : FA port map (A=>sum_0(7), B=>sum_0(6), C_in=>c_out_0(5), S=>sum_1(39) , C_out=>c_out_1(39));
	FA_1_40 : FA port map (A=>pp4(21), B=>pp5(19), C_in=>pp6(17), S=>sum_1(40) , C_out=>c_out_1(40));
	FA_1_41 : FA port map (A=>pp1(27), B=>pp2(25), C_in=>pp3(23), S=>sum_1(41) , C_out=>c_out_1(41));
	FA_1_42 : FA port map (A=>c_out_0(7), B=>c_out_0(6), C_in=>pp0(29), S=>sum_1(42) , C_out=>c_out_1(42));
	FA_1_43 : FA port map (A=>sum_0(10), B=>sum_0(9), C_in=>c_out_0(8), S=>sum_1(43) , C_out=>c_out_1(43));
	FA_1_44 : FA port map (A=>pp3(24), B=>pp4(22), C_in=>pp5(20), S=>sum_1(44) , C_out=>c_out_1(44));
	FA_1_45 : FA port map (A=>pp0(30), B=>pp1(28), C_in=>pp2(26), S=>sum_1(45) , C_out=>c_out_1(45));
	FA_1_46 : FA port map (A=>c_out_0(11), B=>c_out_0(10), C_in=>c_out_0(9), S=>sum_1(46) , C_out=>c_out_1(46));
	FA_1_47 : FA port map (A=>sum_0(14), B=>sum_0(13), C_in=>sum_0(12), S=>sum_1(47) , C_out=>c_out_1(47));
	FA_1_48 : FA port map (A=>pp2(27), B=>pp3(25), C_in=>pp4(23), S=>sum_1(48) , C_out=>c_out_1(48));
	FA_1_49 : FA port map (A=>c_out_0(12), B=>pp0(31), C_in=>pp1(29), S=>sum_1(49) , C_out=>c_out_1(49));
	FA_1_50 : FA port map (A=>c_out_0(15), B=>c_out_0(14), C_in=>c_out_0(13), S=>sum_1(50) , C_out=>c_out_1(50));
	FA_1_51 : FA port map (A=>sum_0(18), B=>sum_0(17), C_in=>sum_0(16), S=>sum_1(51) , C_out=>c_out_1(51));
	FA_1_52 : FA port map (A=>pp2(28), B=>pp3(26), C_in=>pp4(24), S=>sum_1(52) , C_out=>c_out_1(52));
	FA_1_53 : FA port map (A=>c_out_0(16), B=>pp0(32), C_in=>pp1(30), S=>sum_1(53) , C_out=>c_out_1(53));
	FA_1_54 : FA port map (A=>c_out_0(19), B=>c_out_0(18), C_in=>c_out_0(17), S=>sum_1(54) , C_out=>c_out_1(54));
	FA_1_55 : FA port map (A=>sum_0(22), B=>sum_0(21), C_in=>sum_0(20), S=>sum_1(55) , C_out=>c_out_1(55));
	FA_1_56 : FA port map (A=>pp2(29), B=>pp3(27), C_in=>pp4(25), S=>sum_1(56) , C_out=>c_out_1(56));
	FA_1_57 : FA port map (A=>c_out_0(20), B=>s(0), C_in=>pp1(31), S=>sum_1(57) , C_out=>c_out_1(57));
	FA_1_58 : FA port map (A=>c_out_0(23), B=>c_out_0(22), C_in=>c_out_0(21), S=>sum_1(58) , C_out=>c_out_1(58));
	FA_1_59 : FA port map (A=>sum_0(26), B=>sum_0(25), C_in=>sum_0(24), S=>sum_1(59) , C_out=>c_out_1(59));
	FA_1_60 : FA port map (A=>pp2(30), B=>pp3(28), C_in=>pp4(26), S=>sum_1(60) , C_out=>c_out_1(60));
	FA_1_61 : FA port map (A=>c_out_0(24), B=>s(0), C_in=>pp1(32), S=>sum_1(61) , C_out=>c_out_1(61));
	FA_1_62 : FA port map (A=>c_out_0(27), B=>c_out_0(26), C_in=>c_out_0(25), S=>sum_1(62) , C_out=>c_out_1(62));
	FA_1_63 : FA port map (A=>sum_0(30), B=>sum_0(29), C_in=>sum_0(28), S=>sum_1(63) , C_out=>c_out_1(63));
	FA_1_64 : FA port map (A=>pp2(31), B=>pp3(29), C_in=>pp4(27), S=>sum_1(64) , C_out=>c_out_1(64));
	FA_1_65 : FA port map (A=>c_out_0(28), B=>s_n(0), C_in=>s_n(1), S=>sum_1(65) , C_out=>c_out_1(65));
	FA_1_66 : FA port map (A=>c_out_0(31), B=>c_out_0(30), C_in=>c_out_0(29), S=>sum_1(66) , C_out=>c_out_1(66));
	FA_1_67 : FA port map (A=>sum_0(34), B=>sum_0(33), C_in=>sum_0(32), S=>sum_1(67) , C_out=>c_out_1(67));
	FA_1_68 : FA port map (A=>pp3(30), B=>pp4(28), C_in=>pp5(26), S=>sum_1(68) , C_out=>c_out_1(68));
	FA_1_69 : FA port map (A=>c_out_0(32), B=>'1', C_in=>pp2(32), S=>sum_1(69) , C_out=>c_out_1(69));
	FA_1_70 : FA port map (A=>c_out_0(35), B=>c_out_0(34), C_in=>c_out_0(33), S=>sum_1(70) , C_out=>c_out_1(70));
	FA_1_71 : FA port map (A=>sum_0(38), B=>sum_0(37), C_in=>sum_0(36), S=>sum_1(71) , C_out=>c_out_1(71));
	FA_1_72 : FA port map (A=>pp5(27), B=>pp6(25), C_in=>pp7(23), S=>sum_1(72) , C_out=>c_out_1(72));
	FA_1_73 : FA port map (A=>s_n(2), B=>pp3(31), C_in=>pp4(29), S=>sum_1(73) , C_out=>c_out_1(73));
	FA_1_74 : FA port map (A=>c_out_0(38), B=>c_out_0(37), C_in=>c_out_0(36), S=>sum_1(74) , C_out=>c_out_1(74));
	FA_1_75 : FA port map (A=>sum_0(41), B=>sum_0(40), C_in=>c_out_0(39), S=>sum_1(75) , C_out=>c_out_1(75));
	FA_1_76 : FA port map (A=>pp6(26), B=>pp7(24), C_in=>pp8(22), S=>sum_1(76) , C_out=>c_out_1(76));
	FA_1_77 : FA port map (A=>pp3(32), B=>pp4(30), C_in=>pp5(28), S=>sum_1(77) , C_out=>c_out_1(77));
	FA_1_78 : FA port map (A=>c_out_0(41), B=>c_out_0(40), C_in=>'1', S=>sum_1(78) , C_out=>c_out_1(78));
	FA_1_79 : FA port map (A=>sum_0(44), B=>sum_0(43), C_in=>c_out_0(42), S=>sum_1(79) , C_out=>c_out_1(79));
	FA_1_80 : FA port map (A=>pp8(23), B=>pp9(21), C_in=>pp10(19), S=>sum_1(80) , C_out=>c_out_1(80));
	FA_1_81 : FA port map (A=>pp5(29), B=>pp6(27), C_in=>pp7(25), S=>sum_1(81) , C_out=>c_out_1(81));
	FA_1_82 : FA port map (A=>c_out_0(43), B=>s_n(3), C_in=>pp4(31), S=>sum_1(82) , C_out=>c_out_1(82));
	FA_1_83 : FA port map (A=>sum_0(46), B=>c_out_0(45), C_in=>c_out_0(44), S=>sum_1(83) , C_out=>c_out_1(83));
	FA_1_84 : FA port map (A=>pp9(22), B=>pp10(20), C_in=>pp11(18), S=>sum_1(84) , C_out=>c_out_1(84));
	FA_1_85 : FA port map (A=>pp6(28), B=>pp7(26), C_in=>pp8(24), S=>sum_1(85) , C_out=>c_out_1(85));
	FA_1_86 : FA port map (A=>'1', B=>pp4(32), C_in=>pp5(30), S=>sum_1(86) , C_out=>c_out_1(86));
	FA_1_87 : FA port map (A=>sum_0(48), B=>c_out_0(47), C_in=>c_out_0(46), S=>sum_1(87) , C_out=>c_out_1(87));
	FA_1_88 : FA port map (A=>pp11(19), B=>pp12(17), C_in=>pp13(15), S=>sum_1(88) , C_out=>c_out_1(88));
	FA_1_89 : FA port map (A=>pp8(25), B=>pp9(23), C_in=>pp10(21), S=>sum_1(89) , C_out=>c_out_1(89));
	FA_1_90 : FA port map (A=>pp5(31), B=>pp6(29), C_in=>pp7(27), S=>sum_1(90) , C_out=>c_out_1(90));
	FA_1_91 : FA port map (A=>c_out_0(49), B=>c_out_0(48), C_in=>s_n(4), S=>sum_1(91) , C_out=>c_out_1(91));
	FA_1_92 : FA port map (A=>pp12(18), B=>pp13(16), C_in=>pp14(14), S=>sum_1(92) , C_out=>c_out_1(92));
	FA_1_93 : FA port map (A=>pp9(24), B=>pp10(22), C_in=>pp11(20), S=>sum_1(93) , C_out=>c_out_1(93));
	FA_1_94 : FA port map (A=>pp6(30), B=>pp7(28), C_in=>pp8(26), S=>sum_1(94) , C_out=>c_out_1(94));
	FA_1_95 : FA port map (A=>c_out_0(50), B=>'1', C_in=>pp5(32), S=>sum_1(95) , C_out=>c_out_1(95));
	FA_1_96 : FA port map (A=>pp14(15), B=>pp15(13), C_in=>pp16(11), S=>sum_1(96) , C_out=>c_out_1(96));
	FA_1_97 : FA port map (A=>pp11(21), B=>pp12(19), C_in=>pp13(17), S=>sum_1(97) , C_out=>c_out_1(97));
	FA_1_98 : FA port map (A=>pp8(27), B=>pp9(25), C_in=>pp10(23), S=>sum_1(98) , C_out=>c_out_1(98));
	FA_1_99 : FA port map (A=>s_n(5), B=>pp6(31), C_in=>pp7(29), S=>sum_1(99) , C_out=>c_out_1(99));
	FA_1_100 : FA port map (A=>pp14(16), B=>pp15(14), C_in=>pp16(12), S=>sum_1(100) , C_out=>c_out_1(100));
	FA_1_101 : FA port map (A=>pp11(22), B=>pp12(20), C_in=>pp13(18), S=>sum_1(101) , C_out=>c_out_1(101));
	FA_1_102 : FA port map (A=>pp8(28), B=>pp9(26), C_in=>pp10(24), S=>sum_1(102) , C_out=>c_out_1(102));
	HA_1_103 : HA port map (A=>pp6(32), B=>pp7(30), S=>sum_1(103) , C_out=>c_out_1(103));
	FA_1_104 : FA port map (A=>pp14(17), B=>pp15(15), C_in=>pp16(13), S=>sum_1(104) , C_out=>c_out_1(104));
	FA_1_105 : FA port map (A=>pp11(23), B=>pp12(21), C_in=>pp13(19), S=>sum_1(105) , C_out=>c_out_1(105));
	FA_1_106 : FA port map (A=>pp8(29), B=>pp9(27), C_in=>pp10(25), S=>sum_1(106) , C_out=>c_out_1(106));
	FA_1_107 : FA port map (A=>pp14(18), B=>pp15(16), C_in=>pp16(14), S=>sum_1(107) , C_out=>c_out_1(107));
	FA_1_108 : FA port map (A=>pp11(24), B=>pp12(22), C_in=>pp13(20), S=>sum_1(108) , C_out=>c_out_1(108));
	HA_1_109 : HA port map (A=>pp9(28), B=>pp10(26), S=>sum_1(109) , C_out=>c_out_1(109));
	FA_1_110 : FA port map (A=>pp14(19), B=>pp15(17), C_in=>pp16(15), S=>sum_1(110) , C_out=>c_out_1(110));
	FA_1_111 : FA port map (A=>pp11(25), B=>pp12(23), C_in=>pp13(21), S=>sum_1(111) , C_out=>c_out_1(111));
	FA_1_112 : FA port map (A=>pp14(20), B=>pp15(18), C_in=>pp16(16), S=>sum_1(112) , C_out=>c_out_1(112));
	HA_1_113 : HA port map (A=>pp12(24), B=>pp13(22), S=>sum_1(113) , C_out=>c_out_1(113));
	FA_1_114 : FA port map (A=>pp14(21), B=>pp15(19), C_in=>pp16(17), S=>sum_1(114) , C_out=>c_out_1(114));
	HA_1_115 : HA port map (A=>pp15(20), B=>pp16(18), S=>sum_1(115) , C_out=>c_out_1(115));
	HA_2_0 : HA port map (A=>pp5(0), B=>s(5), S=>sum_2(0) , C_out=>c_out_2(0));
	HA_2_1 : HA port map (A=>pp4(3), B=>pp5(1), S=>sum_2(1) , C_out=>c_out_2(1));
	FA_2_2 : FA port map (A=>pp5(2), B=>pp6(0), C_in=>s(6), S=>sum_2(2) , C_out=>c_out_2(2));
	HA_2_3 : HA port map (A=>pp3(6), B=>pp4(4), S=>sum_2(3) , C_out=>c_out_2(3));
	FA_2_4 : FA port map (A=>pp4(5), B=>pp5(3), C_in=>pp6(1), S=>sum_2(4) , C_out=>c_out_2(4));
	HA_2_5 : HA port map (A=>pp2(9), B=>pp3(7), S=>sum_2(5) , C_out=>c_out_2(5));
	FA_2_6 : FA port map (A=>pp6(2), B=>pp7(0), C_in=>s(7), S=>sum_2(6) , C_out=>c_out_2(6));
	FA_2_7 : FA port map (A=>pp3(8), B=>pp4(6), C_in=>pp5(4), S=>sum_2(7) , C_out=>c_out_2(7));
	HA_2_8 : HA port map (A=>pp1(12), B=>pp2(10), S=>sum_2(8) , C_out=>c_out_2(8));
	FA_2_9 : FA port map (A=>pp5(5), B=>pp6(3), C_in=>pp7(1), S=>sum_2(9) , C_out=>c_out_2(9));
	FA_2_10 : FA port map (A=>pp2(11), B=>pp3(9), C_in=>pp4(7), S=>sum_2(10) , C_out=>c_out_2(10));
	HA_2_11 : HA port map (A=>pp0(15), B=>pp1(13), S=>sum_2(11) , C_out=>c_out_2(11));
	FA_2_12 : FA port map (A=>pp5(6), B=>pp6(4), C_in=>pp7(2), S=>sum_2(12) , C_out=>c_out_2(12));
	FA_2_13 : FA port map (A=>pp2(12), B=>pp3(10), C_in=>pp4(8), S=>sum_2(13) , C_out=>c_out_2(13));
	FA_2_14 : FA port map (A=>sum_1(0), B=>pp0(16), C_in=>pp1(14), S=>sum_2(14) , C_out=>c_out_2(14));
	FA_2_15 : FA port map (A=>pp4(9), B=>pp5(7), C_in=>pp6(5), S=>sum_2(15) , C_out=>c_out_2(15));
	FA_2_16 : FA port map (A=>pp1(15), B=>pp2(13), C_in=>pp3(11), S=>sum_2(16) , C_out=>c_out_2(16));
	FA_2_17 : FA port map (A=>sum_1(1), B=>c_out_1(0), C_in=>pp0(17), S=>sum_2(17) , C_out=>c_out_2(17));
	FA_2_18 : FA port map (A=>pp3(12), B=>pp4(10), C_in=>pp5(8), S=>sum_2(18) , C_out=>c_out_2(18));
	FA_2_19 : FA port map (A=>pp0(18), B=>pp1(16), C_in=>pp2(14), S=>sum_2(19) , C_out=>c_out_2(19));
	FA_2_20 : FA port map (A=>sum_1(3), B=>sum_1(2), C_in=>c_out_1(1), S=>sum_2(20) , C_out=>c_out_2(20));
	FA_2_21 : FA port map (A=>pp2(15), B=>pp3(13), C_in=>pp4(11), S=>sum_2(21) , C_out=>c_out_2(21));
	FA_2_22 : FA port map (A=>c_out_1(2), B=>pp0(19), C_in=>pp1(17), S=>sum_2(22) , C_out=>c_out_2(22));
	FA_2_23 : FA port map (A=>sum_1(5), B=>sum_1(4), C_in=>c_out_1(3), S=>sum_2(23) , C_out=>c_out_2(23));
	FA_2_24 : FA port map (A=>pp1(18), B=>pp2(16), C_in=>pp3(14), S=>sum_2(24) , C_out=>c_out_2(24));
	FA_2_25 : FA port map (A=>c_out_1(5), B=>c_out_1(4), C_in=>pp0(20), S=>sum_2(25) , C_out=>c_out_2(25));
	FA_2_26 : FA port map (A=>sum_1(8), B=>sum_1(7), C_in=>sum_1(6), S=>sum_2(26) , C_out=>c_out_2(26));
	FA_2_27 : FA port map (A=>pp0(21), B=>pp1(19), C_in=>pp2(17), S=>sum_2(27) , C_out=>c_out_2(27));
	FA_2_28 : FA port map (A=>c_out_1(8), B=>c_out_1(7), C_in=>c_out_1(6), S=>sum_2(28) , C_out=>c_out_2(28));
	FA_2_29 : FA port map (A=>sum_1(11), B=>sum_1(10), C_in=>sum_1(9), S=>sum_2(29) , C_out=>c_out_2(29));
	FA_2_30 : FA port map (A=>c_out_1(9), B=>pp0(22), C_in=>pp1(20), S=>sum_2(30) , C_out=>c_out_2(30));
	FA_2_31 : FA port map (A=>sum_1(12), B=>c_out_1(11), C_in=>c_out_1(10), S=>sum_2(31) , C_out=>c_out_2(31));
	FA_2_32 : FA port map (A=>sum_1(15), B=>sum_1(14), C_in=>sum_1(13), S=>sum_2(32) , C_out=>c_out_2(32));
	FA_2_33 : FA port map (A=>c_out_1(13), B=>c_out_1(12), C_in=>pp0(23), S=>sum_2(33) , C_out=>c_out_2(33));
	FA_2_34 : FA port map (A=>sum_1(16), B=>c_out_1(15), C_in=>c_out_1(14), S=>sum_2(34) , C_out=>c_out_2(34));
	FA_2_35 : FA port map (A=>sum_1(19), B=>sum_1(18), C_in=>sum_1(17), S=>sum_2(35) , C_out=>c_out_2(35));
	FA_2_36 : FA port map (A=>c_out_1(17), B=>c_out_1(16), C_in=>sum_0(0), S=>sum_2(36) , C_out=>c_out_2(36));
	FA_2_37 : FA port map (A=>sum_1(20), B=>c_out_1(19), C_in=>c_out_1(18), S=>sum_2(37) , C_out=>c_out_2(37));
	FA_2_38 : FA port map (A=>sum_1(23), B=>sum_1(22), C_in=>sum_1(21), S=>sum_2(38) , C_out=>c_out_2(38));
	FA_2_39 : FA port map (A=>c_out_1(21), B=>c_out_1(20), C_in=>sum_0(1), S=>sum_2(39) , C_out=>c_out_2(39));
	FA_2_40 : FA port map (A=>sum_1(24), B=>c_out_1(23), C_in=>c_out_1(22), S=>sum_2(40) , C_out=>c_out_2(40));
	FA_2_41 : FA port map (A=>sum_1(27), B=>sum_1(26), C_in=>sum_1(25), S=>sum_2(41) , C_out=>c_out_2(41));
	FA_2_42 : FA port map (A=>c_out_1(25), B=>c_out_1(24), C_in=>sum_0(3), S=>sum_2(42) , C_out=>c_out_2(42));
	FA_2_43 : FA port map (A=>sum_1(28), B=>c_out_1(27), C_in=>c_out_1(26), S=>sum_2(43) , C_out=>c_out_2(43));
	FA_2_44 : FA port map (A=>sum_1(31), B=>sum_1(30), C_in=>sum_1(29), S=>sum_2(44) , C_out=>c_out_2(44));
	FA_2_45 : FA port map (A=>c_out_1(29), B=>c_out_1(28), C_in=>sum_0(5), S=>sum_2(45) , C_out=>c_out_2(45));
	FA_2_46 : FA port map (A=>sum_1(32), B=>c_out_1(31), C_in=>c_out_1(30), S=>sum_2(46) , C_out=>c_out_2(46));
	FA_2_47 : FA port map (A=>sum_1(35), B=>sum_1(34), C_in=>sum_1(33), S=>sum_2(47) , C_out=>c_out_2(47));
	FA_2_48 : FA port map (A=>c_out_1(33), B=>c_out_1(32), C_in=>sum_0(8), S=>sum_2(48) , C_out=>c_out_2(48));
	FA_2_49 : FA port map (A=>sum_1(36), B=>c_out_1(35), C_in=>c_out_1(34), S=>sum_2(49) , C_out=>c_out_2(49));
	FA_2_50 : FA port map (A=>sum_1(39), B=>sum_1(38), C_in=>sum_1(37), S=>sum_2(50) , C_out=>c_out_2(50));
	FA_2_51 : FA port map (A=>c_out_1(37), B=>c_out_1(36), C_in=>sum_0(11), S=>sum_2(51) , C_out=>c_out_2(51));
	FA_2_52 : FA port map (A=>sum_1(40), B=>c_out_1(39), C_in=>c_out_1(38), S=>sum_2(52) , C_out=>c_out_2(52));
	FA_2_53 : FA port map (A=>sum_1(43), B=>sum_1(42), C_in=>sum_1(41), S=>sum_2(53) , C_out=>c_out_2(53));
	FA_2_54 : FA port map (A=>c_out_1(41), B=>c_out_1(40), C_in=>sum_0(15), S=>sum_2(54) , C_out=>c_out_2(54));
	FA_2_55 : FA port map (A=>sum_1(44), B=>c_out_1(43), C_in=>c_out_1(42), S=>sum_2(55) , C_out=>c_out_2(55));
	FA_2_56 : FA port map (A=>sum_1(47), B=>sum_1(46), C_in=>sum_1(45), S=>sum_2(56) , C_out=>c_out_2(56));
	FA_2_57 : FA port map (A=>c_out_1(45), B=>c_out_1(44), C_in=>sum_0(19), S=>sum_2(57) , C_out=>c_out_2(57));
	FA_2_58 : FA port map (A=>sum_1(48), B=>c_out_1(47), C_in=>c_out_1(46), S=>sum_2(58) , C_out=>c_out_2(58));
	FA_2_59 : FA port map (A=>sum_1(51), B=>sum_1(50), C_in=>sum_1(49), S=>sum_2(59) , C_out=>c_out_2(59));
	FA_2_60 : FA port map (A=>c_out_1(49), B=>c_out_1(48), C_in=>sum_0(23), S=>sum_2(60) , C_out=>c_out_2(60));
	FA_2_61 : FA port map (A=>sum_1(52), B=>c_out_1(51), C_in=>c_out_1(50), S=>sum_2(61) , C_out=>c_out_2(61));
	FA_2_62 : FA port map (A=>sum_1(55), B=>sum_1(54), C_in=>sum_1(53), S=>sum_2(62) , C_out=>c_out_2(62));
	FA_2_63 : FA port map (A=>c_out_1(53), B=>c_out_1(52), C_in=>sum_0(27), S=>sum_2(63) , C_out=>c_out_2(63));
	FA_2_64 : FA port map (A=>sum_1(56), B=>c_out_1(55), C_in=>c_out_1(54), S=>sum_2(64) , C_out=>c_out_2(64));
	FA_2_65 : FA port map (A=>sum_1(59), B=>sum_1(58), C_in=>sum_1(57), S=>sum_2(65) , C_out=>c_out_2(65));
	FA_2_66 : FA port map (A=>c_out_1(57), B=>c_out_1(56), C_in=>sum_0(31), S=>sum_2(66) , C_out=>c_out_2(66));
	FA_2_67 : FA port map (A=>sum_1(60), B=>c_out_1(59), C_in=>c_out_1(58), S=>sum_2(67) , C_out=>c_out_2(67));
	FA_2_68 : FA port map (A=>sum_1(63), B=>sum_1(62), C_in=>sum_1(61), S=>sum_2(68) , C_out=>c_out_2(68));
	FA_2_69 : FA port map (A=>c_out_1(61), B=>c_out_1(60), C_in=>sum_0(35), S=>sum_2(69) , C_out=>c_out_2(69));
	FA_2_70 : FA port map (A=>sum_1(64), B=>c_out_1(63), C_in=>c_out_1(62), S=>sum_2(70) , C_out=>c_out_2(70));
	FA_2_71 : FA port map (A=>sum_1(67), B=>sum_1(66), C_in=>sum_1(65), S=>sum_2(71) , C_out=>c_out_2(71));
	FA_2_72 : FA port map (A=>c_out_1(65), B=>c_out_1(64), C_in=>sum_0(39), S=>sum_2(72) , C_out=>c_out_2(72));
	FA_2_73 : FA port map (A=>sum_1(68), B=>c_out_1(67), C_in=>c_out_1(66), S=>sum_2(73) , C_out=>c_out_2(73));
	FA_2_74 : FA port map (A=>sum_1(71), B=>sum_1(70), C_in=>sum_1(69), S=>sum_2(74) , C_out=>c_out_2(74));
	FA_2_75 : FA port map (A=>c_out_1(69), B=>c_out_1(68), C_in=>sum_0(42), S=>sum_2(75) , C_out=>c_out_2(75));
	FA_2_76 : FA port map (A=>sum_1(72), B=>c_out_1(71), C_in=>c_out_1(70), S=>sum_2(76) , C_out=>c_out_2(76));
	FA_2_77 : FA port map (A=>sum_1(75), B=>sum_1(74), C_in=>sum_1(73), S=>sum_2(77) , C_out=>c_out_2(77));
	FA_2_78 : FA port map (A=>c_out_1(73), B=>c_out_1(72), C_in=>sum_0(45), S=>sum_2(78) , C_out=>c_out_2(78));
	FA_2_79 : FA port map (A=>sum_1(76), B=>c_out_1(75), C_in=>c_out_1(74), S=>sum_2(79) , C_out=>c_out_2(79));
	FA_2_80 : FA port map (A=>sum_1(79), B=>sum_1(78), C_in=>sum_1(77), S=>sum_2(80) , C_out=>c_out_2(80));
	FA_2_81 : FA port map (A=>c_out_1(77), B=>c_out_1(76), C_in=>sum_0(47), S=>sum_2(81) , C_out=>c_out_2(81));
	FA_2_82 : FA port map (A=>sum_1(80), B=>c_out_1(79), C_in=>c_out_1(78), S=>sum_2(82) , C_out=>c_out_2(82));
	FA_2_83 : FA port map (A=>sum_1(83), B=>sum_1(82), C_in=>sum_1(81), S=>sum_2(83) , C_out=>c_out_2(83));
	FA_2_84 : FA port map (A=>c_out_1(81), B=>c_out_1(80), C_in=>sum_0(49), S=>sum_2(84) , C_out=>c_out_2(84));
	FA_2_85 : FA port map (A=>sum_1(84), B=>c_out_1(83), C_in=>c_out_1(82), S=>sum_2(85) , C_out=>c_out_2(85));
	FA_2_86 : FA port map (A=>sum_1(87), B=>sum_1(86), C_in=>sum_1(85), S=>sum_2(86) , C_out=>c_out_2(86));
	FA_2_87 : FA port map (A=>c_out_1(85), B=>c_out_1(84), C_in=>sum_0(50), S=>sum_2(87) , C_out=>c_out_2(87));
	FA_2_88 : FA port map (A=>sum_1(88), B=>c_out_1(87), C_in=>c_out_1(86), S=>sum_2(88) , C_out=>c_out_2(88));
	FA_2_89 : FA port map (A=>sum_1(91), B=>sum_1(90), C_in=>sum_1(89), S=>sum_2(89) , C_out=>c_out_2(89));
	FA_2_90 : FA port map (A=>c_out_1(89), B=>c_out_1(88), C_in=>sum_0(51), S=>sum_2(90) , C_out=>c_out_2(90));
	FA_2_91 : FA port map (A=>sum_1(92), B=>c_out_1(91), C_in=>c_out_1(90), S=>sum_2(91) , C_out=>c_out_2(91));
	FA_2_92 : FA port map (A=>sum_1(95), B=>sum_1(94), C_in=>sum_1(93), S=>sum_2(92) , C_out=>c_out_2(92));
	FA_2_93 : FA port map (A=>c_out_1(93), B=>c_out_1(92), C_in=>c_out_0(51), S=>sum_2(93) , C_out=>c_out_2(93));
	FA_2_94 : FA port map (A=>sum_1(96), B=>c_out_1(95), C_in=>c_out_1(94), S=>sum_2(94) , C_out=>c_out_2(94));
	FA_2_95 : FA port map (A=>sum_1(99), B=>sum_1(98), C_in=>sum_1(97), S=>sum_2(95) , C_out=>c_out_2(95));
	FA_2_96 : FA port map (A=>c_out_1(97), B=>c_out_1(96), C_in=>'1', S=>sum_2(96) , C_out=>c_out_2(96));
	FA_2_97 : FA port map (A=>sum_1(100), B=>c_out_1(99), C_in=>c_out_1(98), S=>sum_2(97) , C_out=>c_out_2(97));
	FA_2_98 : FA port map (A=>sum_1(103), B=>sum_1(102), C_in=>sum_1(101), S=>sum_2(98) , C_out=>c_out_2(98));
	FA_2_99 : FA port map (A=>c_out_1(100), B=>s_n(6), C_in=>pp7(31), S=>sum_2(99) , C_out=>c_out_2(99));
	FA_2_100 : FA port map (A=>c_out_1(103), B=>c_out_1(102), C_in=>c_out_1(101), S=>sum_2(100) , C_out=>c_out_2(100));
	FA_2_101 : FA port map (A=>sum_1(106), B=>sum_1(105), C_in=>sum_1(104), S=>sum_2(101) , C_out=>c_out_2(101));
	FA_2_102 : FA port map (A=>'1', B=>pp7(32), C_in=>pp8(30), S=>sum_2(102) , C_out=>c_out_2(102));
	FA_2_103 : FA port map (A=>c_out_1(106), B=>c_out_1(105), C_in=>c_out_1(104), S=>sum_2(103) , C_out=>c_out_2(103));
	FA_2_104 : FA port map (A=>sum_1(109), B=>sum_1(108), C_in=>sum_1(107), S=>sum_2(104) , C_out=>c_out_2(104));
	FA_2_105 : FA port map (A=>pp8(31), B=>pp9(29), C_in=>pp10(27), S=>sum_2(105) , C_out=>c_out_2(105));
	FA_2_106 : FA port map (A=>c_out_1(108), B=>c_out_1(107), C_in=>s_n(7), S=>sum_2(106) , C_out=>c_out_2(106));
	FA_2_107 : FA port map (A=>sum_1(111), B=>sum_1(110), C_in=>c_out_1(109), S=>sum_2(107) , C_out=>c_out_2(107));
	FA_2_108 : FA port map (A=>pp9(30), B=>pp10(28), C_in=>pp11(26), S=>sum_2(108) , C_out=>c_out_2(108));
	FA_2_109 : FA port map (A=>c_out_1(110), B=>'1', C_in=>pp8(32), S=>sum_2(109) , C_out=>c_out_2(109));
	FA_2_110 : FA port map (A=>sum_1(113), B=>sum_1(112), C_in=>c_out_1(111), S=>sum_2(110) , C_out=>c_out_2(110));
	FA_2_111 : FA port map (A=>pp11(27), B=>pp12(25), C_in=>pp13(23), S=>sum_2(111) , C_out=>c_out_2(111));
	FA_2_112 : FA port map (A=>s_n(8), B=>pp9(31), C_in=>pp10(29), S=>sum_2(112) , C_out=>c_out_2(112));
	FA_2_113 : FA port map (A=>sum_1(114), B=>c_out_1(113), C_in=>c_out_1(112), S=>sum_2(113) , C_out=>c_out_2(113));
	FA_2_114 : FA port map (A=>pp12(26), B=>pp13(24), C_in=>pp14(22), S=>sum_2(114) , C_out=>c_out_2(114));
	FA_2_115 : FA port map (A=>pp9(32), B=>pp10(30), C_in=>pp11(28), S=>sum_2(115) , C_out=>c_out_2(115));
	FA_2_116 : FA port map (A=>sum_1(115), B=>c_out_1(114), C_in=>'1', S=>sum_2(116) , C_out=>c_out_2(116));
	FA_2_117 : FA port map (A=>pp14(23), B=>pp15(21), C_in=>pp16(19), S=>sum_2(117) , C_out=>c_out_2(117));
	FA_2_118 : FA port map (A=>pp11(29), B=>pp12(27), C_in=>pp13(25), S=>sum_2(118) , C_out=>c_out_2(118));
	FA_2_119 : FA port map (A=>c_out_1(115), B=>s_n(9), C_in=>pp10(31), S=>sum_2(119) , C_out=>c_out_2(119));
	FA_2_120 : FA port map (A=>pp14(24), B=>pp15(22), C_in=>pp16(20), S=>sum_2(120) , C_out=>c_out_2(120));
	FA_2_121 : FA port map (A=>pp11(30), B=>pp12(28), C_in=>pp13(26), S=>sum_2(121) , C_out=>c_out_2(121));
	HA_2_122 : HA port map (A=>'1', B=>pp10(32), S=>sum_2(122) , C_out=>c_out_2(122));
	FA_2_123 : FA port map (A=>pp14(25), B=>pp15(23), C_in=>pp16(21), S=>sum_2(123) , C_out=>c_out_2(123));
	FA_2_124 : FA port map (A=>pp11(31), B=>pp12(29), C_in=>pp13(27), S=>sum_2(124) , C_out=>c_out_2(124));
	FA_2_125 : FA port map (A=>pp14(26), B=>pp15(24), C_in=>pp16(22), S=>sum_2(125) , C_out=>c_out_2(125));
	HA_2_126 : HA port map (A=>pp12(30), B=>pp13(28), S=>sum_2(126) , C_out=>c_out_2(126));
	FA_2_127 : FA port map (A=>pp14(27), B=>pp15(25), C_in=>pp16(23), S=>sum_2(127) , C_out=>c_out_2(127));
	HA_2_128 : HA port map (A=>pp15(26), B=>pp16(24), S=>sum_2(128) , C_out=>c_out_2(128));
	HA_3_0 : HA port map (A=>pp3(0), B=>s(3), S=>sum_3(0) , C_out=>c_out_3(0));
	HA_3_1 : HA port map (A=>pp2(3), B=>pp3(1), S=>sum_3(1) , C_out=>c_out_3(1));
	FA_3_2 : FA port map (A=>pp3(2), B=>pp4(0), C_in=>s(4), S=>sum_3(2) , C_out=>c_out_3(2));
	HA_3_3 : HA port map (A=>pp1(6), B=>pp2(4), S=>sum_3(3) , C_out=>c_out_3(3));
	FA_3_4 : FA port map (A=>pp2(5), B=>pp3(3), C_in=>pp4(1), S=>sum_3(4) , C_out=>c_out_3(4));
	HA_3_5 : HA port map (A=>pp0(9), B=>pp1(7), S=>sum_3(5) , C_out=>c_out_3(5));
	FA_3_6 : FA port map (A=>pp2(6), B=>pp3(4), C_in=>pp4(2), S=>sum_3(6) , C_out=>c_out_3(6));
	FA_3_7 : FA port map (A=>sum_2(0), B=>pp0(10), C_in=>pp1(8), S=>sum_3(7) , C_out=>c_out_3(7));
	FA_3_8 : FA port map (A=>pp1(9), B=>pp2(7), C_in=>pp3(5), S=>sum_3(8) , C_out=>c_out_3(8));
	FA_3_9 : FA port map (A=>sum_2(1), B=>c_out_2(0), C_in=>pp0(11), S=>sum_3(9) , C_out=>c_out_3(9));
	FA_3_10 : FA port map (A=>pp0(12), B=>pp1(10), C_in=>pp2(8), S=>sum_3(10) , C_out=>c_out_3(10));
	FA_3_11 : FA port map (A=>sum_2(3), B=>sum_2(2), C_in=>c_out_2(1), S=>sum_3(11) , C_out=>c_out_3(11));
	FA_3_12 : FA port map (A=>c_out_2(2), B=>pp0(13), C_in=>pp1(11), S=>sum_3(12) , C_out=>c_out_3(12));
	FA_3_13 : FA port map (A=>sum_2(5), B=>sum_2(4), C_in=>c_out_2(3), S=>sum_3(13) , C_out=>c_out_3(13));
	FA_3_14 : FA port map (A=>c_out_2(5), B=>c_out_2(4), C_in=>pp0(14), S=>sum_3(14) , C_out=>c_out_3(14));
	FA_3_15 : FA port map (A=>sum_2(8), B=>sum_2(7), C_in=>sum_2(6), S=>sum_3(15) , C_out=>c_out_3(15));
	FA_3_16 : FA port map (A=>c_out_2(8), B=>c_out_2(7), C_in=>c_out_2(6), S=>sum_3(16) , C_out=>c_out_3(16));
	FA_3_17 : FA port map (A=>sum_2(11), B=>sum_2(10), C_in=>sum_2(9), S=>sum_3(17) , C_out=>c_out_3(17));
	FA_3_18 : FA port map (A=>c_out_2(11), B=>c_out_2(10), C_in=>c_out_2(9), S=>sum_3(18) , C_out=>c_out_3(18));
	FA_3_19 : FA port map (A=>sum_2(14), B=>sum_2(13), C_in=>sum_2(12), S=>sum_3(19) , C_out=>c_out_3(19));
	FA_3_20 : FA port map (A=>c_out_2(14), B=>c_out_2(13), C_in=>c_out_2(12), S=>sum_3(20) , C_out=>c_out_3(20));
	FA_3_21 : FA port map (A=>sum_2(17), B=>sum_2(16), C_in=>sum_2(15), S=>sum_3(21) , C_out=>c_out_3(21));
	FA_3_22 : FA port map (A=>c_out_2(17), B=>c_out_2(16), C_in=>c_out_2(15), S=>sum_3(22) , C_out=>c_out_3(22));
	FA_3_23 : FA port map (A=>sum_2(20), B=>sum_2(19), C_in=>sum_2(18), S=>sum_3(23) , C_out=>c_out_3(23));
	FA_3_24 : FA port map (A=>c_out_2(20), B=>c_out_2(19), C_in=>c_out_2(18), S=>sum_3(24) , C_out=>c_out_3(24));
	FA_3_25 : FA port map (A=>sum_2(23), B=>sum_2(22), C_in=>sum_2(21), S=>sum_3(25) , C_out=>c_out_3(25));
	FA_3_26 : FA port map (A=>c_out_2(23), B=>c_out_2(22), C_in=>c_out_2(21), S=>sum_3(26) , C_out=>c_out_3(26));
	FA_3_27 : FA port map (A=>sum_2(26), B=>sum_2(25), C_in=>sum_2(24), S=>sum_3(27) , C_out=>c_out_3(27));
	FA_3_28 : FA port map (A=>c_out_2(26), B=>c_out_2(25), C_in=>c_out_2(24), S=>sum_3(28) , C_out=>c_out_3(28));
	FA_3_29 : FA port map (A=>sum_2(29), B=>sum_2(28), C_in=>sum_2(27), S=>sum_3(29) , C_out=>c_out_3(29));
	FA_3_30 : FA port map (A=>c_out_2(29), B=>c_out_2(28), C_in=>c_out_2(27), S=>sum_3(30) , C_out=>c_out_3(30));
	FA_3_31 : FA port map (A=>sum_2(32), B=>sum_2(31), C_in=>sum_2(30), S=>sum_3(31) , C_out=>c_out_3(31));
	FA_3_32 : FA port map (A=>c_out_2(32), B=>c_out_2(31), C_in=>c_out_2(30), S=>sum_3(32) , C_out=>c_out_3(32));
	FA_3_33 : FA port map (A=>sum_2(35), B=>sum_2(34), C_in=>sum_2(33), S=>sum_3(33) , C_out=>c_out_3(33));
	FA_3_34 : FA port map (A=>c_out_2(35), B=>c_out_2(34), C_in=>c_out_2(33), S=>sum_3(34) , C_out=>c_out_3(34));
	FA_3_35 : FA port map (A=>sum_2(38), B=>sum_2(37), C_in=>sum_2(36), S=>sum_3(35) , C_out=>c_out_3(35));
	FA_3_36 : FA port map (A=>c_out_2(38), B=>c_out_2(37), C_in=>c_out_2(36), S=>sum_3(36) , C_out=>c_out_3(36));
	FA_3_37 : FA port map (A=>sum_2(41), B=>sum_2(40), C_in=>sum_2(39), S=>sum_3(37) , C_out=>c_out_3(37));
	FA_3_38 : FA port map (A=>c_out_2(41), B=>c_out_2(40), C_in=>c_out_2(39), S=>sum_3(38) , C_out=>c_out_3(38));
	FA_3_39 : FA port map (A=>sum_2(44), B=>sum_2(43), C_in=>sum_2(42), S=>sum_3(39) , C_out=>c_out_3(39));
	FA_3_40 : FA port map (A=>c_out_2(44), B=>c_out_2(43), C_in=>c_out_2(42), S=>sum_3(40) , C_out=>c_out_3(40));
	FA_3_41 : FA port map (A=>sum_2(47), B=>sum_2(46), C_in=>sum_2(45), S=>sum_3(41) , C_out=>c_out_3(41));
	FA_3_42 : FA port map (A=>c_out_2(47), B=>c_out_2(46), C_in=>c_out_2(45), S=>sum_3(42) , C_out=>c_out_3(42));
	FA_3_43 : FA port map (A=>sum_2(50), B=>sum_2(49), C_in=>sum_2(48), S=>sum_3(43) , C_out=>c_out_3(43));
	FA_3_44 : FA port map (A=>c_out_2(50), B=>c_out_2(49), C_in=>c_out_2(48), S=>sum_3(44) , C_out=>c_out_3(44));
	FA_3_45 : FA port map (A=>sum_2(53), B=>sum_2(52), C_in=>sum_2(51), S=>sum_3(45) , C_out=>c_out_3(45));
	FA_3_46 : FA port map (A=>c_out_2(53), B=>c_out_2(52), C_in=>c_out_2(51), S=>sum_3(46) , C_out=>c_out_3(46));
	FA_3_47 : FA port map (A=>sum_2(56), B=>sum_2(55), C_in=>sum_2(54), S=>sum_3(47) , C_out=>c_out_3(47));
	FA_3_48 : FA port map (A=>c_out_2(56), B=>c_out_2(55), C_in=>c_out_2(54), S=>sum_3(48) , C_out=>c_out_3(48));
	FA_3_49 : FA port map (A=>sum_2(59), B=>sum_2(58), C_in=>sum_2(57), S=>sum_3(49) , C_out=>c_out_3(49));
	FA_3_50 : FA port map (A=>c_out_2(59), B=>c_out_2(58), C_in=>c_out_2(57), S=>sum_3(50) , C_out=>c_out_3(50));
	FA_3_51 : FA port map (A=>sum_2(62), B=>sum_2(61), C_in=>sum_2(60), S=>sum_3(51) , C_out=>c_out_3(51));
	FA_3_52 : FA port map (A=>c_out_2(62), B=>c_out_2(61), C_in=>c_out_2(60), S=>sum_3(52) , C_out=>c_out_3(52));
	FA_3_53 : FA port map (A=>sum_2(65), B=>sum_2(64), C_in=>sum_2(63), S=>sum_3(53) , C_out=>c_out_3(53));
	FA_3_54 : FA port map (A=>c_out_2(65), B=>c_out_2(64), C_in=>c_out_2(63), S=>sum_3(54) , C_out=>c_out_3(54));
	FA_3_55 : FA port map (A=>sum_2(68), B=>sum_2(67), C_in=>sum_2(66), S=>sum_3(55) , C_out=>c_out_3(55));
	FA_3_56 : FA port map (A=>c_out_2(68), B=>c_out_2(67), C_in=>c_out_2(66), S=>sum_3(56) , C_out=>c_out_3(56));
	FA_3_57 : FA port map (A=>sum_2(71), B=>sum_2(70), C_in=>sum_2(69), S=>sum_3(57) , C_out=>c_out_3(57));
	FA_3_58 : FA port map (A=>c_out_2(71), B=>c_out_2(70), C_in=>c_out_2(69), S=>sum_3(58) , C_out=>c_out_3(58));
	FA_3_59 : FA port map (A=>sum_2(74), B=>sum_2(73), C_in=>sum_2(72), S=>sum_3(59) , C_out=>c_out_3(59));
	FA_3_60 : FA port map (A=>c_out_2(74), B=>c_out_2(73), C_in=>c_out_2(72), S=>sum_3(60) , C_out=>c_out_3(60));
	FA_3_61 : FA port map (A=>sum_2(77), B=>sum_2(76), C_in=>sum_2(75), S=>sum_3(61) , C_out=>c_out_3(61));
	FA_3_62 : FA port map (A=>c_out_2(77), B=>c_out_2(76), C_in=>c_out_2(75), S=>sum_3(62) , C_out=>c_out_3(62));
	FA_3_63 : FA port map (A=>sum_2(80), B=>sum_2(79), C_in=>sum_2(78), S=>sum_3(63) , C_out=>c_out_3(63));
	FA_3_64 : FA port map (A=>c_out_2(80), B=>c_out_2(79), C_in=>c_out_2(78), S=>sum_3(64) , C_out=>c_out_3(64));
	FA_3_65 : FA port map (A=>sum_2(83), B=>sum_2(82), C_in=>sum_2(81), S=>sum_3(65) , C_out=>c_out_3(65));
	FA_3_66 : FA port map (A=>c_out_2(83), B=>c_out_2(82), C_in=>c_out_2(81), S=>sum_3(66) , C_out=>c_out_3(66));
	FA_3_67 : FA port map (A=>sum_2(86), B=>sum_2(85), C_in=>sum_2(84), S=>sum_3(67) , C_out=>c_out_3(67));
	FA_3_68 : FA port map (A=>c_out_2(86), B=>c_out_2(85), C_in=>c_out_2(84), S=>sum_3(68) , C_out=>c_out_3(68));
	FA_3_69 : FA port map (A=>sum_2(89), B=>sum_2(88), C_in=>sum_2(87), S=>sum_3(69) , C_out=>c_out_3(69));
	FA_3_70 : FA port map (A=>c_out_2(89), B=>c_out_2(88), C_in=>c_out_2(87), S=>sum_3(70) , C_out=>c_out_3(70));
	FA_3_71 : FA port map (A=>sum_2(92), B=>sum_2(91), C_in=>sum_2(90), S=>sum_3(71) , C_out=>c_out_3(71));
	FA_3_72 : FA port map (A=>c_out_2(92), B=>c_out_2(91), C_in=>c_out_2(90), S=>sum_3(72) , C_out=>c_out_3(72));
	FA_3_73 : FA port map (A=>sum_2(95), B=>sum_2(94), C_in=>sum_2(93), S=>sum_3(73) , C_out=>c_out_3(73));
	FA_3_74 : FA port map (A=>c_out_2(95), B=>c_out_2(94), C_in=>c_out_2(93), S=>sum_3(74) , C_out=>c_out_3(74));
	FA_3_75 : FA port map (A=>sum_2(98), B=>sum_2(97), C_in=>sum_2(96), S=>sum_3(75) , C_out=>c_out_3(75));
	FA_3_76 : FA port map (A=>c_out_2(98), B=>c_out_2(97), C_in=>c_out_2(96), S=>sum_3(76) , C_out=>c_out_3(76));
	FA_3_77 : FA port map (A=>sum_2(101), B=>sum_2(100), C_in=>sum_2(99), S=>sum_3(77) , C_out=>c_out_3(77));
	FA_3_78 : FA port map (A=>c_out_2(101), B=>c_out_2(100), C_in=>c_out_2(99), S=>sum_3(78) , C_out=>c_out_3(78));
	FA_3_79 : FA port map (A=>sum_2(104), B=>sum_2(103), C_in=>sum_2(102), S=>sum_3(79) , C_out=>c_out_3(79));
	FA_3_80 : FA port map (A=>c_out_2(104), B=>c_out_2(103), C_in=>c_out_2(102), S=>sum_3(80) , C_out=>c_out_3(80));
	FA_3_81 : FA port map (A=>sum_2(107), B=>sum_2(106), C_in=>sum_2(105), S=>sum_3(81) , C_out=>c_out_3(81));
	FA_3_82 : FA port map (A=>c_out_2(107), B=>c_out_2(106), C_in=>c_out_2(105), S=>sum_3(82) , C_out=>c_out_3(82));
	FA_3_83 : FA port map (A=>sum_2(110), B=>sum_2(109), C_in=>sum_2(108), S=>sum_3(83) , C_out=>c_out_3(83));
	FA_3_84 : FA port map (A=>c_out_2(110), B=>c_out_2(109), C_in=>c_out_2(108), S=>sum_3(84) , C_out=>c_out_3(84));
	FA_3_85 : FA port map (A=>sum_2(113), B=>sum_2(112), C_in=>sum_2(111), S=>sum_3(85) , C_out=>c_out_3(85));
	FA_3_86 : FA port map (A=>c_out_2(113), B=>c_out_2(112), C_in=>c_out_2(111), S=>sum_3(86) , C_out=>c_out_3(86));
	FA_3_87 : FA port map (A=>sum_2(116), B=>sum_2(115), C_in=>sum_2(114), S=>sum_3(87) , C_out=>c_out_3(87));
	FA_3_88 : FA port map (A=>c_out_2(116), B=>c_out_2(115), C_in=>c_out_2(114), S=>sum_3(88) , C_out=>c_out_3(88));
	FA_3_89 : FA port map (A=>sum_2(119), B=>sum_2(118), C_in=>sum_2(117), S=>sum_3(89) , C_out=>c_out_3(89));
	FA_3_90 : FA port map (A=>c_out_2(119), B=>c_out_2(118), C_in=>c_out_2(117), S=>sum_3(90) , C_out=>c_out_3(90));
	FA_3_91 : FA port map (A=>sum_2(122), B=>sum_2(121), C_in=>sum_2(120), S=>sum_3(91) , C_out=>c_out_3(91));
	FA_3_92 : FA port map (A=>c_out_2(121), B=>c_out_2(120), C_in=>s_n(10), S=>sum_3(92) , C_out=>c_out_3(92));
	FA_3_93 : FA port map (A=>sum_2(124), B=>sum_2(123), C_in=>c_out_2(122), S=>sum_3(93) , C_out=>c_out_3(93));
	FA_3_94 : FA port map (A=>c_out_2(123), B=>'1', C_in=>pp11(32), S=>sum_3(94) , C_out=>c_out_3(94));
	FA_3_95 : FA port map (A=>sum_2(126), B=>sum_2(125), C_in=>c_out_2(124), S=>sum_3(95) , C_out=>c_out_3(95));
	FA_3_96 : FA port map (A=>s_n(11), B=>pp12(31), C_in=>pp13(29), S=>sum_3(96) , C_out=>c_out_3(96));
	FA_3_97 : FA port map (A=>sum_2(127), B=>c_out_2(126), C_in=>c_out_2(125), S=>sum_3(97) , C_out=>c_out_3(97));
	FA_3_98 : FA port map (A=>pp12(32), B=>pp13(30), C_in=>pp14(28), S=>sum_3(98) , C_out=>c_out_3(98));
	FA_3_99 : FA port map (A=>sum_2(128), B=>c_out_2(127), C_in=>'1', S=>sum_3(99) , C_out=>c_out_3(99));
	FA_3_100 : FA port map (A=>pp14(29), B=>pp15(27), C_in=>pp16(25), S=>sum_3(100) , C_out=>c_out_3(100));
	FA_3_101 : FA port map (A=>c_out_2(128), B=>s_n(12), C_in=>pp13(31), S=>sum_3(101) , C_out=>c_out_3(101));
	FA_3_102 : FA port map (A=>pp14(30), B=>pp15(28), C_in=>pp16(26), S=>sum_3(102) , C_out=>c_out_3(102));
	HA_3_103 : HA port map (A=>'1', B=>pp13(32), S=>sum_3(103) , C_out=>c_out_3(103));
	FA_3_104 : FA port map (A=>pp14(31), B=>pp15(29), C_in=>pp16(27), S=>sum_3(104) , C_out=>c_out_3(104));
	HA_3_105 : HA port map (A=>pp15(30), B=>pp16(28), S=>sum_3(105) , C_out=>c_out_3(105));
	HA_4_0 : HA port map (A=>pp2(0), B=>s(2), S=>sum_4(0) , C_out=>c_out_4(0));
	HA_4_1 : HA port map (A=>pp1(3), B=>pp2(1), S=>sum_4(1) , C_out=>c_out_4(1));
	FA_4_2 : FA port map (A=>pp0(6), B=>pp1(4), C_in=>pp2(2), S=>sum_4(2) , C_out=>c_out_4(2));
	FA_4_3 : FA port map (A=>c_out_3(0), B=>pp0(7), C_in=>pp1(5), S=>sum_4(3) , C_out=>c_out_4(3));
	FA_4_4 : FA port map (A=>sum_3(2), B=>c_out_3(1), C_in=>pp0(8), S=>sum_4(4) , C_out=>c_out_4(4));
	FA_4_5 : FA port map (A=>sum_3(4), B=>c_out_3(3), C_in=>c_out_3(2), S=>sum_4(5) , C_out=>c_out_4(5));
	FA_4_6 : FA port map (A=>sum_3(6), B=>c_out_3(5), C_in=>c_out_3(4), S=>sum_4(6) , C_out=>c_out_4(6));
	FA_4_7 : FA port map (A=>sum_3(8), B=>c_out_3(7), C_in=>c_out_3(6), S=>sum_4(7) , C_out=>c_out_4(7));
	FA_4_8 : FA port map (A=>sum_3(10), B=>c_out_3(9), C_in=>c_out_3(8), S=>sum_4(8) , C_out=>c_out_4(8));
	FA_4_9 : FA port map (A=>sum_3(12), B=>c_out_3(11), C_in=>c_out_3(10), S=>sum_4(9) , C_out=>c_out_4(9));
	FA_4_10 : FA port map (A=>sum_3(14), B=>c_out_3(13), C_in=>c_out_3(12), S=>sum_4(10) , C_out=>c_out_4(10));
	FA_4_11 : FA port map (A=>sum_3(16), B=>c_out_3(15), C_in=>c_out_3(14), S=>sum_4(11) , C_out=>c_out_4(11));
	FA_4_12 : FA port map (A=>sum_3(18), B=>c_out_3(17), C_in=>c_out_3(16), S=>sum_4(12) , C_out=>c_out_4(12));
	FA_4_13 : FA port map (A=>sum_3(20), B=>c_out_3(19), C_in=>c_out_3(18), S=>sum_4(13) , C_out=>c_out_4(13));
	FA_4_14 : FA port map (A=>sum_3(22), B=>c_out_3(21), C_in=>c_out_3(20), S=>sum_4(14) , C_out=>c_out_4(14));
	FA_4_15 : FA port map (A=>sum_3(24), B=>c_out_3(23), C_in=>c_out_3(22), S=>sum_4(15) , C_out=>c_out_4(15));
	FA_4_16 : FA port map (A=>sum_3(26), B=>c_out_3(25), C_in=>c_out_3(24), S=>sum_4(16) , C_out=>c_out_4(16));
	FA_4_17 : FA port map (A=>sum_3(28), B=>c_out_3(27), C_in=>c_out_3(26), S=>sum_4(17) , C_out=>c_out_4(17));
	FA_4_18 : FA port map (A=>sum_3(30), B=>c_out_3(29), C_in=>c_out_3(28), S=>sum_4(18) , C_out=>c_out_4(18));
	FA_4_19 : FA port map (A=>sum_3(32), B=>c_out_3(31), C_in=>c_out_3(30), S=>sum_4(19) , C_out=>c_out_4(19));
	FA_4_20 : FA port map (A=>sum_3(34), B=>c_out_3(33), C_in=>c_out_3(32), S=>sum_4(20) , C_out=>c_out_4(20));
	FA_4_21 : FA port map (A=>sum_3(36), B=>c_out_3(35), C_in=>c_out_3(34), S=>sum_4(21) , C_out=>c_out_4(21));
	FA_4_22 : FA port map (A=>sum_3(38), B=>c_out_3(37), C_in=>c_out_3(36), S=>sum_4(22) , C_out=>c_out_4(22));
	FA_4_23 : FA port map (A=>sum_3(40), B=>c_out_3(39), C_in=>c_out_3(38), S=>sum_4(23) , C_out=>c_out_4(23));
	FA_4_24 : FA port map (A=>sum_3(42), B=>c_out_3(41), C_in=>c_out_3(40), S=>sum_4(24) , C_out=>c_out_4(24));
	FA_4_25 : FA port map (A=>sum_3(44), B=>c_out_3(43), C_in=>c_out_3(42), S=>sum_4(25) , C_out=>c_out_4(25));
	FA_4_26 : FA port map (A=>sum_3(46), B=>c_out_3(45), C_in=>c_out_3(44), S=>sum_4(26) , C_out=>c_out_4(26));
	FA_4_27 : FA port map (A=>sum_3(48), B=>c_out_3(47), C_in=>c_out_3(46), S=>sum_4(27) , C_out=>c_out_4(27));
	FA_4_28 : FA port map (A=>sum_3(50), B=>c_out_3(49), C_in=>c_out_3(48), S=>sum_4(28) , C_out=>c_out_4(28));
	FA_4_29 : FA port map (A=>sum_3(52), B=>c_out_3(51), C_in=>c_out_3(50), S=>sum_4(29) , C_out=>c_out_4(29));
	FA_4_30 : FA port map (A=>sum_3(54), B=>c_out_3(53), C_in=>c_out_3(52), S=>sum_4(30) , C_out=>c_out_4(30));
	FA_4_31 : FA port map (A=>sum_3(56), B=>c_out_3(55), C_in=>c_out_3(54), S=>sum_4(31) , C_out=>c_out_4(31));
	FA_4_32 : FA port map (A=>sum_3(58), B=>c_out_3(57), C_in=>c_out_3(56), S=>sum_4(32) , C_out=>c_out_4(32));
	FA_4_33 : FA port map (A=>sum_3(60), B=>c_out_3(59), C_in=>c_out_3(58), S=>sum_4(33) , C_out=>c_out_4(33));
	FA_4_34 : FA port map (A=>sum_3(62), B=>c_out_3(61), C_in=>c_out_3(60), S=>sum_4(34) , C_out=>c_out_4(34));
	FA_4_35 : FA port map (A=>sum_3(64), B=>c_out_3(63), C_in=>c_out_3(62), S=>sum_4(35) , C_out=>c_out_4(35));
	FA_4_36 : FA port map (A=>sum_3(66), B=>c_out_3(65), C_in=>c_out_3(64), S=>sum_4(36) , C_out=>c_out_4(36));
	FA_4_37 : FA port map (A=>sum_3(68), B=>c_out_3(67), C_in=>c_out_3(66), S=>sum_4(37) , C_out=>c_out_4(37));
	FA_4_38 : FA port map (A=>sum_3(70), B=>c_out_3(69), C_in=>c_out_3(68), S=>sum_4(38) , C_out=>c_out_4(38));
	FA_4_39 : FA port map (A=>sum_3(72), B=>c_out_3(71), C_in=>c_out_3(70), S=>sum_4(39) , C_out=>c_out_4(39));
	FA_4_40 : FA port map (A=>sum_3(74), B=>c_out_3(73), C_in=>c_out_3(72), S=>sum_4(40) , C_out=>c_out_4(40));
	FA_4_41 : FA port map (A=>sum_3(76), B=>c_out_3(75), C_in=>c_out_3(74), S=>sum_4(41) , C_out=>c_out_4(41));
	FA_4_42 : FA port map (A=>sum_3(78), B=>c_out_3(77), C_in=>c_out_3(76), S=>sum_4(42) , C_out=>c_out_4(42));
	FA_4_43 : FA port map (A=>sum_3(80), B=>c_out_3(79), C_in=>c_out_3(78), S=>sum_4(43) , C_out=>c_out_4(43));
	FA_4_44 : FA port map (A=>sum_3(82), B=>c_out_3(81), C_in=>c_out_3(80), S=>sum_4(44) , C_out=>c_out_4(44));
	FA_4_45 : FA port map (A=>sum_3(84), B=>c_out_3(83), C_in=>c_out_3(82), S=>sum_4(45) , C_out=>c_out_4(45));
	FA_4_46 : FA port map (A=>sum_3(86), B=>c_out_3(85), C_in=>c_out_3(84), S=>sum_4(46) , C_out=>c_out_4(46));
	FA_4_47 : FA port map (A=>sum_3(88), B=>c_out_3(87), C_in=>c_out_3(86), S=>sum_4(47) , C_out=>c_out_4(47));
	FA_4_48 : FA port map (A=>sum_3(90), B=>c_out_3(89), C_in=>c_out_3(88), S=>sum_4(48) , C_out=>c_out_4(48));
	FA_4_49 : FA port map (A=>sum_3(92), B=>c_out_3(91), C_in=>c_out_3(90), S=>sum_4(49) , C_out=>c_out_4(49));
	FA_4_50 : FA port map (A=>sum_3(94), B=>c_out_3(93), C_in=>c_out_3(92), S=>sum_4(50) , C_out=>c_out_4(50));
	FA_4_51 : FA port map (A=>sum_3(96), B=>c_out_3(95), C_in=>c_out_3(94), S=>sum_4(51) , C_out=>c_out_4(51));
	FA_4_52 : FA port map (A=>sum_3(98), B=>c_out_3(97), C_in=>c_out_3(96), S=>sum_4(52) , C_out=>c_out_4(52));
	FA_4_53 : FA port map (A=>sum_3(100), B=>c_out_3(99), C_in=>c_out_3(98), S=>sum_4(53) , C_out=>c_out_4(53));
	FA_4_54 : FA port map (A=>sum_3(102), B=>c_out_3(101), C_in=>c_out_3(100), S=>sum_4(54) , C_out=>c_out_4(54));
	FA_4_55 : FA port map (A=>c_out_3(103), B=>c_out_3(102), C_in=>s_n(13), S=>sum_4(55) , C_out=>c_out_4(55));
	FA_4_56 : FA port map (A=>c_out_3(104), B=>'1', C_in=>pp14(32), S=>sum_4(56) , C_out=>c_out_4(56));
	FA_4_57 : FA port map (A=>s_n(14), B=>pp15(31), C_in=>pp16(29), S=>sum_4(57) , C_out=>c_out_4(57));
	HA_4_58 : HA port map (A=>pp15(32), B=>pp16(30), S=>sum_4(58) , C_out=>c_out_4(58));
	HA_5_0 : HA port map (A=>pp1(0), B=>s(1), S=>sum_5(0) , C_out=>c_out_5(0));
	HA_5_1 : HA port map (A=>pp0(3), B=>pp1(1), S=>sum_5(1) , C_out=>c_out_5(1));
	FA_5_2 : FA port map (A=>sum_4(0), B=>pp0(4), C_in=>pp1(2), S=>sum_5(2) , C_out=>c_out_5(2));
	FA_5_3 : FA port map (A=>sum_4(1), B=>c_out_4(0), C_in=>pp0(5), S=>sum_5(3) , C_out=>c_out_5(3));
	FA_5_4 : FA port map (A=>sum_4(2), B=>c_out_4(1), C_in=>sum_3(0), S=>sum_5(4) , C_out=>c_out_5(4));
	FA_5_5 : FA port map (A=>sum_4(3), B=>c_out_4(2), C_in=>sum_3(1), S=>sum_5(5) , C_out=>c_out_5(5));
	FA_5_6 : FA port map (A=>sum_4(4), B=>c_out_4(3), C_in=>sum_3(3), S=>sum_5(6) , C_out=>c_out_5(6));
	FA_5_7 : FA port map (A=>sum_4(5), B=>c_out_4(4), C_in=>sum_3(5), S=>sum_5(7) , C_out=>c_out_5(7));
	FA_5_8 : FA port map (A=>sum_4(6), B=>c_out_4(5), C_in=>sum_3(7), S=>sum_5(8) , C_out=>c_out_5(8));
	FA_5_9 : FA port map (A=>sum_4(7), B=>c_out_4(6), C_in=>sum_3(9), S=>sum_5(9) , C_out=>c_out_5(9));
	FA_5_10 : FA port map (A=>sum_4(8), B=>c_out_4(7), C_in=>sum_3(11), S=>sum_5(10) , C_out=>c_out_5(10));
	FA_5_11 : FA port map (A=>sum_4(9), B=>c_out_4(8), C_in=>sum_3(13), S=>sum_5(11) , C_out=>c_out_5(11));
	FA_5_12 : FA port map (A=>sum_4(10), B=>c_out_4(9), C_in=>sum_3(15), S=>sum_5(12) , C_out=>c_out_5(12));
	FA_5_13 : FA port map (A=>sum_4(11), B=>c_out_4(10), C_in=>sum_3(17), S=>sum_5(13) , C_out=>c_out_5(13));
	FA_5_14 : FA port map (A=>sum_4(12), B=>c_out_4(11), C_in=>sum_3(19), S=>sum_5(14) , C_out=>c_out_5(14));
	FA_5_15 : FA port map (A=>sum_4(13), B=>c_out_4(12), C_in=>sum_3(21), S=>sum_5(15) , C_out=>c_out_5(15));
	FA_5_16 : FA port map (A=>sum_4(14), B=>c_out_4(13), C_in=>sum_3(23), S=>sum_5(16) , C_out=>c_out_5(16));
	FA_5_17 : FA port map (A=>sum_4(15), B=>c_out_4(14), C_in=>sum_3(25), S=>sum_5(17) , C_out=>c_out_5(17));
	FA_5_18 : FA port map (A=>sum_4(16), B=>c_out_4(15), C_in=>sum_3(27), S=>sum_5(18) , C_out=>c_out_5(18));
	FA_5_19 : FA port map (A=>sum_4(17), B=>c_out_4(16), C_in=>sum_3(29), S=>sum_5(19) , C_out=>c_out_5(19));
	FA_5_20 : FA port map (A=>sum_4(18), B=>c_out_4(17), C_in=>sum_3(31), S=>sum_5(20) , C_out=>c_out_5(20));
	FA_5_21 : FA port map (A=>sum_4(19), B=>c_out_4(18), C_in=>sum_3(33), S=>sum_5(21) , C_out=>c_out_5(21));
	FA_5_22 : FA port map (A=>sum_4(20), B=>c_out_4(19), C_in=>sum_3(35), S=>sum_5(22) , C_out=>c_out_5(22));
	FA_5_23 : FA port map (A=>sum_4(21), B=>c_out_4(20), C_in=>sum_3(37), S=>sum_5(23) , C_out=>c_out_5(23));
	FA_5_24 : FA port map (A=>sum_4(22), B=>c_out_4(21), C_in=>sum_3(39), S=>sum_5(24) , C_out=>c_out_5(24));
	FA_5_25 : FA port map (A=>sum_4(23), B=>c_out_4(22), C_in=>sum_3(41), S=>sum_5(25) , C_out=>c_out_5(25));
	FA_5_26 : FA port map (A=>sum_4(24), B=>c_out_4(23), C_in=>sum_3(43), S=>sum_5(26) , C_out=>c_out_5(26));
	FA_5_27 : FA port map (A=>sum_4(25), B=>c_out_4(24), C_in=>sum_3(45), S=>sum_5(27) , C_out=>c_out_5(27));
	FA_5_28 : FA port map (A=>sum_4(26), B=>c_out_4(25), C_in=>sum_3(47), S=>sum_5(28) , C_out=>c_out_5(28));
	FA_5_29 : FA port map (A=>sum_4(27), B=>c_out_4(26), C_in=>sum_3(49), S=>sum_5(29) , C_out=>c_out_5(29));
	FA_5_30 : FA port map (A=>sum_4(28), B=>c_out_4(27), C_in=>sum_3(51), S=>sum_5(30) , C_out=>c_out_5(30));
	FA_5_31 : FA port map (A=>sum_4(29), B=>c_out_4(28), C_in=>sum_3(53), S=>sum_5(31) , C_out=>c_out_5(31));
	FA_5_32 : FA port map (A=>sum_4(30), B=>c_out_4(29), C_in=>sum_3(55), S=>sum_5(32) , C_out=>c_out_5(32));
	FA_5_33 : FA port map (A=>sum_4(31), B=>c_out_4(30), C_in=>sum_3(57), S=>sum_5(33) , C_out=>c_out_5(33));
	FA_5_34 : FA port map (A=>sum_4(32), B=>c_out_4(31), C_in=>sum_3(59), S=>sum_5(34) , C_out=>c_out_5(34));
	FA_5_35 : FA port map (A=>sum_4(33), B=>c_out_4(32), C_in=>sum_3(61), S=>sum_5(35) , C_out=>c_out_5(35));
	FA_5_36 : FA port map (A=>sum_4(34), B=>c_out_4(33), C_in=>sum_3(63), S=>sum_5(36) , C_out=>c_out_5(36));
	FA_5_37 : FA port map (A=>sum_4(35), B=>c_out_4(34), C_in=>sum_3(65), S=>sum_5(37) , C_out=>c_out_5(37));
	FA_5_38 : FA port map (A=>sum_4(36), B=>c_out_4(35), C_in=>sum_3(67), S=>sum_5(38) , C_out=>c_out_5(38));
	FA_5_39 : FA port map (A=>sum_4(37), B=>c_out_4(36), C_in=>sum_3(69), S=>sum_5(39) , C_out=>c_out_5(39));
	FA_5_40 : FA port map (A=>sum_4(38), B=>c_out_4(37), C_in=>sum_3(71), S=>sum_5(40) , C_out=>c_out_5(40));
	FA_5_41 : FA port map (A=>sum_4(39), B=>c_out_4(38), C_in=>sum_3(73), S=>sum_5(41) , C_out=>c_out_5(41));
	FA_5_42 : FA port map (A=>sum_4(40), B=>c_out_4(39), C_in=>sum_3(75), S=>sum_5(42) , C_out=>c_out_5(42));
	FA_5_43 : FA port map (A=>sum_4(41), B=>c_out_4(40), C_in=>sum_3(77), S=>sum_5(43) , C_out=>c_out_5(43));
	FA_5_44 : FA port map (A=>sum_4(42), B=>c_out_4(41), C_in=>sum_3(79), S=>sum_5(44) , C_out=>c_out_5(44));
	FA_5_45 : FA port map (A=>sum_4(43), B=>c_out_4(42), C_in=>sum_3(81), S=>sum_5(45) , C_out=>c_out_5(45));
	FA_5_46 : FA port map (A=>sum_4(44), B=>c_out_4(43), C_in=>sum_3(83), S=>sum_5(46) , C_out=>c_out_5(46));
	FA_5_47 : FA port map (A=>sum_4(45), B=>c_out_4(44), C_in=>sum_3(85), S=>sum_5(47) , C_out=>c_out_5(47));
	FA_5_48 : FA port map (A=>sum_4(46), B=>c_out_4(45), C_in=>sum_3(87), S=>sum_5(48) , C_out=>c_out_5(48));
	FA_5_49 : FA port map (A=>sum_4(47), B=>c_out_4(46), C_in=>sum_3(89), S=>sum_5(49) , C_out=>c_out_5(49));
	FA_5_50 : FA port map (A=>sum_4(48), B=>c_out_4(47), C_in=>sum_3(91), S=>sum_5(50) , C_out=>c_out_5(50));
	FA_5_51 : FA port map (A=>sum_4(49), B=>c_out_4(48), C_in=>sum_3(93), S=>sum_5(51) , C_out=>c_out_5(51));
	FA_5_52 : FA port map (A=>sum_4(50), B=>c_out_4(49), C_in=>sum_3(95), S=>sum_5(52) , C_out=>c_out_5(52));
	FA_5_53 : FA port map (A=>sum_4(51), B=>c_out_4(50), C_in=>sum_3(97), S=>sum_5(53) , C_out=>c_out_5(53));
	FA_5_54 : FA port map (A=>sum_4(52), B=>c_out_4(51), C_in=>sum_3(99), S=>sum_5(54) , C_out=>c_out_5(54));
	FA_5_55 : FA port map (A=>sum_4(53), B=>c_out_4(52), C_in=>sum_3(101), S=>sum_5(55) , C_out=>c_out_5(55));
	FA_5_56 : FA port map (A=>sum_4(54), B=>c_out_4(53), C_in=>sum_3(103), S=>sum_5(56) , C_out=>c_out_5(56));
	FA_5_57 : FA port map (A=>sum_4(55), B=>c_out_4(54), C_in=>sum_3(104), S=>sum_5(57) , C_out=>c_out_5(57));
	FA_5_58 : FA port map (A=>sum_4(56), B=>c_out_4(55), C_in=>sum_3(105), S=>sum_5(58) , C_out=>c_out_5(58));
	FA_5_59 : FA port map (A=>sum_4(57), B=>c_out_4(56), C_in=>c_out_3(105), S=>sum_5(59) , C_out=>c_out_5(59));
	FA_5_60 : FA port map (A=>sum_4(58), B=>c_out_4(57), C_in=>'1', S=>sum_5(60) , C_out=>c_out_5(60));
	FA_5_61 : FA port map (A=>c_out_4(58), B=>s_n(15), C_in=>pp16(31), S=>sum_5(61) , C_out=>c_out_5(61));

	HA_6 : HA port map (A=>pp0(0), B=>s(0), S=>sum_6, C_out=>c_out_6);

	addend1_out <= sum_5(61) & sum_5(60) & sum_5(59) & sum_5(58) & sum_5(57) & sum_5(56) & sum_5(55) & sum_5(54) & sum_5(53) & sum_5(52) & sum_5(51) & sum_5(50) & sum_5(49) & sum_5(48) & sum_5(47) & sum_5(46) & sum_5(45) & sum_5(44) & sum_5(43) & sum_5(42) & sum_5(41) & sum_5(40) & sum_5(39) & sum_5(38) & sum_5(37) & sum_5(36) & sum_5(35) & sum_5(34) & sum_5(33) & sum_5(32) & sum_5(31) & sum_5(30) & sum_5(29) & sum_5(28) & sum_5(27) & sum_5(26) & sum_5(25) & sum_5(24) & sum_5(23) & sum_5(22) & sum_5(21) & sum_5(20) & sum_5(19) & sum_5(18) & sum_5(17) & sum_5(16) & sum_5(15) & sum_5(14) & sum_5(13) & sum_5(12) & sum_5(11) & sum_5(10) & sum_5(9) & sum_5(8) & sum_5(7) & sum_5(6) & sum_5(5) & sum_5(4) & sum_5(3) & sum_5(2) & sum_5(1) & sum_5(0) & c_out_6;

	addend2_out <= c_out_5(60) & c_out_5(59) & c_out_5(58) & c_out_5(57) & c_out_5(56) & c_out_5(55) & c_out_5(54) & c_out_5(53) & c_out_5(52) & c_out_5(51) & c_out_5(50) & c_out_5(49) & c_out_5(48) & c_out_5(47) & c_out_5(46) & c_out_5(45) & c_out_5(44) & c_out_5(43) & c_out_5(42) & c_out_5(41) & c_out_5(40) & c_out_5(39) & c_out_5(38) & c_out_5(37) & c_out_5(36) & c_out_5(35) & c_out_5(34) & c_out_5(33) & c_out_5(32) & c_out_5(31) & c_out_5(30) & c_out_5(29) & c_out_5(28) & c_out_5(27) & c_out_5(26) & c_out_5(25) & c_out_5(24) & c_out_5(23) & c_out_5(22) & c_out_5(21) & c_out_5(20) & c_out_5(19) & c_out_5(18) & c_out_5(17) & c_out_5(16) & c_out_5(15) & c_out_5(14) & c_out_5(13) & c_out_5(12) & c_out_5(11) & c_out_5(10) & c_out_5(9) & c_out_5(8) & c_out_5(7) & c_out_5(6) & c_out_5(5) & c_out_5(4) & c_out_5(3) & c_out_5(2) & c_out_5(1) & c_out_5(0) & pp0(2) & pp0(1);

	M_lsb <= sum_6;

END struct;