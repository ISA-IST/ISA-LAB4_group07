class packet_in extends uvm_sequence_item;
    rand integer unsigned A;
    rand integer unsigned B;

//	constraint my_A { A > 0 ;}
//	constraint my_B { B > 0 ;}

    `uvm_object_utils_begin(packet_in)
        `uvm_field_int(A, UVM_ALL_ON|UVM_HEX)
        `uvm_field_int(B, UVM_ALL_ON|UVM_HEX)
    `uvm_object_utils_end

    function new(string name="packet_in");
        super.new(name);
    endfunction: new
endclass: packet_in
